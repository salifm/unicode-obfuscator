// Copyright 2020 Salif Mehmed
// Licensed under the EUPL

module unicode_obfuscator

const (
	chars_map = [
		['a', 'а'], ['c', 'с'], ['e', 'е'], ['k', 'к'], ['n', 'п'],
		['o', 'о'], ['p', 'р'], ['x', 'х'], ['y', 'у'], ['A', 'А'],
		['C', 'С'], ['E', 'Е'], ['H', 'Н'], ['K', 'К'], ['O', 'О'],
		['P', 'Р'], ['T', 'Т'], ['X', 'Х'], ['Y', 'У']
	]
)
