// Copyright 2020 Salif Mehmed
// Licensed under the EUPL

module unicode_obfuscator

const (
	invisible_char = "​"
	invisible_char_code = 8203
)
