module main

fn main() {
	println("under construction")
	exit(1)
}
