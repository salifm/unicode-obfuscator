// Copyright 2020 Salif Mehmed
// Licensed under the EUPL

module unicode_obfuscator

pub fn parse_args(args []string) []string {
	r := args
	return r
}

pub fn exec_args(args []string) int {
	println("under construction")
	return 1
}
